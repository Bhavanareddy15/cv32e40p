`ifndef ALU_PKG_SV
`define ALU_PKG_SV

package alu_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import cv32e40p_pkg::*;

  `include "alu_seq_item.sv"
  `include "alu_config.sv"
  `include "alu_sequencer.sv"
  `include "alu_sequences.sv"
  `include "alu_driver.sv"
  `include "alu_monitor.sv"
  `include "alu_agent.sv"
  `include "alu_env.sv"
  `include "alu_test.sv"

endpackage

`endif
